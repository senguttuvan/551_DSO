
module cmd_module(clk,rst_n,SPI_done,cmd,cmd_rdy,SPI_data,ss,wrt_SPI,EEP_data,send_resp,clr_cmd_rdy,resp_sent,resp_to_send,
                  trig_cfg,trig_pos,decimator_reg,capture_done,ch1_rdata,ch2_rdata,ch3_rdata,addr,trace_end,
									clr_capture_done,dump_en);

input clk,rst_n,SPI_done;
input cmd_rdy;
input [23:0] cmd;
input resp_sent;
input [7:0] EEP_data;
input capture_done;                               // set trig_cfg[5] to 0 , whenever capture_done is asserted
input [8:0] trace_end;
input [7:0] ch1_rdata,ch2_rdata,ch3_rdata;

output reg [8:0] trig_pos;                       //inputs to the capture module
output reg [3:0] decimator_reg;
output reg [7:0] trig_cfg;
output reg [7:0] resp_to_send;                   //flopped version of resp_data
output [15:0] SPI_data;
output [2:0] ss;
output wrt_SPI,send_resp;
output clr_cmd_rdy;
output reg [8:0] addr;
output reg clr_capture_done,dump_en;

   //////////////////////////////////////////////////////////////////////////
  // Interconnects between modules...declare any wire types you need here //
 //////////////////////////////////////////////////////////////////////////

 reg set_dec,cfg_pot,set_trig_cfg,set_pos, set_sum,set_prod;												//control signals 
 reg capture_ch1_gain, capture_ch2_gain,capture_ch3_gain;         //control signals for gain of the channels
 reg [15:0] SPI_data;	
 reg [2:0] ss;
 reg wrt_SPI,send_resp,SPI_done_ff;                                                 
 reg clr_cmd_rdy;
 reg [2:0] ch1_gain,ch2_gain,ch3_gain;
 reg [7:0] offset,gain, resp_data;
 reg flop_offset,flop_gain, flop_resp;
 wire [7:0] raw , adder_out;																			// Output/Input to offset correction module                                             
 wire [7:0] corrected;
 reg strt_addrcnt,en_addrcnt,set_channel;
 reg [1:0] chnl;                                                  //to store cc ie channel 
 reg capture_done_ff;                                           
 reg [7:0] sum;
 reg [7:0] prod;

 localparam DUMP_CHN 		= 4'h1;
 localparam CFG_GAIN 		= 4'h2;
 localparam SET_TRIG 		= 4'h3;
 localparam CFG_TRG_POS = 4'h4;
 localparam SET_DEC 		= 4'h5;
 localparam WRITE_TRIG 	= 4'h6;
 localparam READ_TRIG 	= 4'h7;
 localparam WRT_EEP  		= 4'h8;
 localparam RD_EEP   		= 4'h9;

 typedef enum reg [3:0] {CMD_DISPATCH,RD_OFFSET1,RD_GAIN1,RD_OFFSET2,DUMP1,DUMP2,DUMP3,CFG_GAIN2,SET_TRIG2,WRT_EEP2,RD_EEP2,RD_EEP3} state_t;

 state_t state,nstate;


////////////////////////////////////
///////ACK and NACK params/////////
localparam ACK = 8'hA5;
localparam NACK = 8'hEE;
//////////////////////////////////

   /////////////////////////////////////////////
  // Instantiation of gain correction logic  //
 /////////////////////////////////////////////

 assign raw =  (~cmd[9] & ~cmd[8]) ? ch1_rdata : 
								(~cmd[9] & cmd[8]) ?  ch2_rdata : ch3_rdata;

// calib_eep icorr(.raw(raw),.off(offset),.gain(gain),.corrected(corrected));
 saturation_adder iadd(.raw(raw),.off(offset) ,.sums(adder_out));
 saturation_multiplier imul(.sums(sum), .gain(gain) ,.corrected(corrected));

  ///////////////////////////////////
  // Logic for Command processing //
  /////////////////////////////////


 always_ff @(posedge clk, negedge rst_n)
		if (!rst_n)
			sum <= 0;
		else if(set_sum)
			sum <= adder_out;

always_ff @ (posedge clk,negedge rst_n)                 
	if (!rst_n)
		clr_capture_done <= 0;
 else if(set_trig_cfg)
		clr_capture_done <= ~cmd[13];
 else
		clr_capture_done <= 0;

always_ff @ (posedge clk,negedge rst_n)                 
	if (!rst_n)
		SPI_done_ff <= 0;
 else 
		SPI_done_ff	<= SPI_done;




// resp data is flopped as resp_to_send

 always_ff @(posedge clk, negedge rst_n) 
    if(~rst_n)
      resp_to_send <= 8'h00;
    else if(flop_resp)
      resp_to_send <= resp_data;

///////////////////////////////////////////////////////////////////																			
///////////////////////address ofthe EEPROM///////////////////////
///////////////////////////////////////////////////////////////////

	always_ff @(posedge clk, negedge rst_n) 
		if(~rst_n)
			addr <= 9'h000;
		else if(strt_addrcnt)
			addr <= trace_end + 1;
		else if(en_addrcnt)
			addr <= addr + 1;

///////////////////////////////////////////////////////////////////
/////////////////////Decimator Register///////////////////////////
//////////////////////////////////////////////////////////////////	

always_ff @ (posedge clk,negedge rst_n)
	if (!rst_n)
		decimator_reg <= 4'b0000;
	else if(set_dec)
		decimator_reg <= cmd[3:0];

///////////////////////////////////////////////////////////////////
///////////////////////////trigger position register///////////////
////////////////////////////////////////////////////////////////////
always_ff @ (posedge clk,negedge rst_n)
	if (!rst_n)
		trig_pos <= 9'h000;
	else if(set_pos)
		trig_pos <= cmd[8:0];

////////////////////////////////////////////////////////////////////////
/////////////////////Trigger configure register during write/////////
//////////////////////////////////////////////////////////////////////
always_ff @ (posedge clk,negedge rst_n)                 
	if (!rst_n)
		trig_cfg <= 6'h00;
 else if(set_trig_cfg)
		trig_cfg[5:0]	<= cmd[13:8];     
  else if( capture_done )
		trig_cfg[5] <= 1;
	else if( ~capture_done )
		trig_cfg[5] <= 0;

/////////////////////////////////////////////////////////////////////////
//////////////////Implementation of state machine///////////////////////
////////////////////////////////////////////////////////////////////////
always_ff @ (posedge clk,negedge rst_n)
	if (!rst_n)
		state <= CMD_DISPATCH;
	else
		state <= nstate;

///////////////////////////////////////////////////////////////////
/////////////////////Gain of channel 1////////////////////////////
//////////////////////////////////////////////////////////////////
always_ff @ (posedge clk,negedge rst_n)
	if (!rst_n)
		ch1_gain <= 3'b000;
	else if(capture_ch1_gain)
		ch1_gain <= cmd[12:10];

/////////////////////////////////////////////////////////////////
//////////////////Gain of channel 2////////////////////////////
//////////////////////////////////////////////////////////////
always_ff @ (posedge clk,negedge rst_n)
	if (!rst_n)
		ch2_gain <= 3'b000;
	else if(capture_ch2_gain)
		ch2_gain <= cmd[12:10];

//////////////////////////////////////////////////////////////////
//////////////////Gain of channel 3////////////////////////////
//////////////////////////////////////////////////////////////
always_ff @ (posedge clk,negedge rst_n)
	if (!rst_n)
		ch3_gain <= 3'b000;
	else if(capture_ch3_gain)
		ch3_gain <= cmd[12:10];

////////////////////////////////////////////////////////////////
//////////////////Offset from calibration EEPROM///////////////
//////////////////////////////////////////////////////////////
always_ff @ (posedge clk,negedge rst_n)
	if (!rst_n)
		offset <= 8'h00;
	else if(flop_offset)
		offset <= EEP_data;

//////////////////////////////////////////////////////////////
//////////////////Gain from calibration EEPROM///////////////
////////////////////////////////////////////////////////////
always_ff @ (posedge clk,negedge rst_n)
	if (!rst_n)
		gain <= 8'h00;
	else if(flop_gain)
		gain <= EEP_data;


/////////////////////////////////////////////////
//////////////////channel ie cc ///////////////
//////////////////////////////////////////////
/*always_ff @ (posedge clk,negedge rst_n)
	if (!rst_n)
		chnl <= 2'b00;
	else if(set_channel)
		chnl <= cmd[9:8];
*/

/////////////////////////////////////////////////////
//////////////////Combinational block///////////////
///////////////////////////////////////////////////
always_comb 
begin	

 SPI_data = 16'h0000;                      //Default values
 ss = 3'b000;
 wrt_SPI = 0;
 flop_resp = 0;
 send_resp = 0;
 clr_cmd_rdy = 0;
 resp_data = 8'hA5;
 capture_ch1_gain = 0;
 capture_ch2_gain = 0;
 capture_ch3_gain = 0;
 flop_offset = 0;
 flop_gain = 0;
 strt_addrcnt = 0;
 en_addrcnt = 0;
 set_channel = 0;
 set_dec=0;
 set_trig_cfg=0;
 set_pos=0;
 dump_en = 0;
 set_sum = 0;
 set_prod = 0;

case (state)
			CMD_DISPATCH : begin                                      //if state is CMD_DISPATCH check for cmd_rdy
											if (cmd_rdy) begin												//if cmd_rdy is high check the first byte of cmd
												case (cmd[19:16])

														DUMP_CHN : begin
																								 wrt_SPI = 1;            //set channel used for assigning cc (ie channel) in chnl
																								 ss = 3'b100;
																								 set_channel = 1;
																	case (cmd[9:8])
																				2'b00 : begin
																								SPI_data = {4'h0,ch1_gain,1'b0,8'h00};          
																								end
																				2'b01 : begin
																								SPI_data = {4'h1,ch2_gain,1'b0,8'h00};		
																								end
																				2'b10 : begin
																								SPI_data = {4'h2,ch3_gain,1'b0,8'h00};		
																								end
																	endcase
															nstate = RD_OFFSET1;                                     //go to offset state 
															end

															CFG_GAIN : begin
																									wrt_SPI = 1;
																									///// ss is determined from cmd[9:8]//////////////////////////////////////
                                                  ////and the gain for each channel is obtained from cmd using control signal 
                                                  ////capture_ch_gain////////////////////////////////////////////////////////
																	case (cmd[9:8])         
																				2'b00 : begin
																								ss = 3'b001;
																								capture_ch1_gain = 1;
																								end
																				2'b01 : begin
																								ss = 3'b010;
																								capture_ch2_gain  = 1;
																								end
																				default : begin                               
																								ss = 3'b011;
																								capture_ch3_gain  = 1;	            
																								end
																	endcase
			
																							////// SPI data to send based on ggg bits/////////////////
																	case (cmd[12:10])
																				3'b000 : SPI_data = 16'h1302;
																				3'b001 : SPI_data = 16'h1305;
																				3'b010 : SPI_data = 16'h1309;
																				3'b011 : SPI_data = 16'h1314;
																				3'b100 : SPI_data = 16'h1328;
																				3'b101 : SPI_data = 16'h1346;
																				3'b110 : SPI_data = 16'h136B;
																				3'b111 : SPI_data = 16'h13DD;
																endcase
						
															nstate = CFG_GAIN2;            
				  															end
																				
						
			 											SET_TRIG : begin                                              ///////trigger level is set///////////
																			ss = 3'b000;
																			SPI_data = {8'h13,cmd[7:0]};                      /////data is sent on the SPI bus///////
        	 														wrt_SPI = 1;
																			nstate = SET_TRIG2;
				  														end
				
																
                            CFG_TRG_POS:begin
																				set_pos=1;              ///when set_pos is high a positive ACK is sent//////
            														resp_data = ACK;      
            														flop_resp = 1;          ////flop resp is used to flop resp_data////////
            														send_resp = 1;          ////send _resp goes high/////////
            														clr_cmd_rdy = 1;
																				nstate=CMD_DISPATCH;     //////at the end clr_cmd_rdy goes high/////////
																				end

														SET_DEC:		begin
																				set_dec=1;                ////////same as CFG_TRG_POS////////////////
            														resp_data = ACK; 
            														flop_resp = 1;
            														send_resp = 1;
            														clr_cmd_rdy = 1;
																				nstate=CMD_DISPATCH;
																				end

														WRITE_TRIG: begin
																				set_trig_cfg=1;								////when set_trig_cfg goes high the trig_cfg is written///////
              													resp_data = ACK;
              													flop_resp = 1;
              													send_resp = 1;
              													clr_cmd_rdy = 1;
																				nstate=CMD_DISPATCH;
																				end

														READ_TRIG:	begin                                                    ///trig_cfg is read////////////////////////
																			resp_data=trig_cfg;  
            													flop_resp = 1;                     
																			send_resp=1;
           													 	clr_cmd_rdy = 1;
																			nstate=CMD_DISPATCH;
																			end	

														WRT_EEP : begin
					 														wrt_SPI = 1;
																			ss = 3'b100;			                                 // select EEPROM on SPI bus
																			SPI_data = {2'b01,cmd[13:0]};	                    // addresss is in 13:8 , data to write is in 7:0
																			nstate = WRT_EEP2;
				   														end

			  										RD_EEP : 	begin
					 														wrt_SPI = 1;
																			ss = 3'b100;			                               // select EEPROM on SPI bus
																			SPI_data = {2'b00,cmd[13:0]};	                  // addresss is in 13:8 
																			nstate = RD_EEP2;
				  														end

			  									  default : begin	                                            // unkown command so neg ack
																		resp_data = NACK;
            												flop_resp = 1;
            												send_resp = 1;
            												clr_cmd_rdy = 1;
																		ss = 3'b000;
																		capture_ch1_gain = 0;
																		capture_ch2_gain = 0;
																		capture_ch3_gain = 0;
																		SPI_data = 16'h0000;
																		wrt_SPI = 0;
																		nstate = CMD_DISPATCH;
			  														end
												endcase
										end
						else 
												nstate = CMD_DISPATCH;
		
					end


///////////////////////////////////////////
/////   read offset command is sent  /////
/////////////////////////////////////////


					RD_OFFSET1 :  begin
											 if (SPI_done_ff && SPI_done) begin                                //SPI sends out junk value so goes to next state ie RD_GAIN1 when SPI_done is high
													 nstate = RD_GAIN1;	
													 wrt_SPI = 1;		
		 	 										 ss = 3'b100;
														case (cmd[9:8])                             //data is written on the SPI bus
																	2'b00 : begin
																					SPI_data = {4'h0,ch1_gain,1'b1,8'h00};
																					end
																	2'b01 : begin
																					SPI_data = {4'h1,ch2_gain,1'b1,8'h00};						
																					end
																	2'b10 : begin
																					SPI_data = {4'h2,ch3_gain,1'b1,8'h00};						
																					end
														endcase
									  		  end else begin
				 									 ss = 3'b100;	                                                 // select EEPROM on SPI bus
													 nstate = RD_OFFSET1;                          //otherwise stays in same state///////////////////
											 end
	 										 end


/////////////////////////////////////////////////////////////////////
/////  Offset value is read and the read gain command is sent  /////
///////////////////////////////////////////////////////////////////


 				 RD_GAIN1 : 	begin
											if (SPI_done_ff && SPI_done) begin
												nstate = RD_OFFSET2;                        //SPI sends the offset value that is obtained when flop_offset is high////
												flop_gain = 1;                            ///then goes to next state ie OFFSET2
												wrt_SPI = 1;
												ss = 3'b100;	
 												SPI_data = 16'h0000;               //junk value is sent to SPI
											end
											else begin
												nstate = RD_GAIN1;
												ss = 3'b100;
											end
	 										end


////////////////////////////////////////////////////////////////
///////////  Wait state till the gain value is read  //////////
//////////////////////////////////////////////////////////////



					RD_OFFSET2 : begin                                        //SPI sends the gain value and it is stored when flop_gain is high
											if(SPI_done_ff && SPI_done) begin
																	nstate = DUMP1;
																	flop_offset = 1;
																	dump_en = 1;
		  														strt_addrcnt = 1;             //addr is assigned to trace_end + 1 
													end
											else begin
															ss = 3'b100;	                  	// select EEPROM on SPI bus
															nstate = RD_OFFSET2;
													end
											end




//////////////////////////////////////////////////////////////////////////////////////////////////////////
/////////////if addr is equal to trace, dumping is over and clr_capture_done bit goes high///////////
////////////////////////////////////////////////////////////////////////////////////////////////////////


					DUMP1 : begin
									dump_en = 1;
									if(addr == trace_end) begin             
      																clr_cmd_rdy = 1;
																			nstate = CMD_DISPATCH;
   																			end
									else begin																			//otherwise the corrected value is sent out the UART and it goes to DUMP3
														nstate = DUMP2;
														set_sum = 1;
//		  																send_resp = 1;
												end
									 	end

					DUMP2 : begin
											dump_en = 1;
											nstate = DUMP3;
											resp_data = corrected;
	   									flop_resp = 1;
											send_resp = 1;
									end


/////////////////////////////////////////////////////////////////////////////////////////////////////////////
/////////////////////if UART sends the resp_sent signal then the process continues until addr equals trace_end///
////////////////////At each stage addr is incremented///////////////////////////////////////////////////////

  				DUMP3 : begin
									dump_en = 1;
											if(resp_sent) begin
			 													nstate = DUMP1;
			 													en_addrcnt = 1;
																			end
	 										else
			 													nstate = DUMP3;
									end


//////////////////////////////////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////wait state for configure gain state///////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////
					CFG_GAIN2 : begin
											   if(SPI_done) begin
        													 clr_cmd_rdy = 1;
        													 resp_data = ACK;
        													 flop_resp = 1;
		    													 send_resp = 1;
																	 nstate = CMD_DISPATCH;
    															    end
											   else  begin
																		ss = (~cmd[9] & ~cmd[8]) ? 3'b001 : 
																				 ((~cmd[9] & cmd[8]) ?  3'b010 : 3'b011 );
	     															nstate = CFG_GAIN2;
															end
											end

////////////////////////////////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////wait state for set trigger level////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////////////////////
 					SET_TRIG2 : begin
												 if(SPI_done) begin
        													clr_cmd_rdy = 1;
        													resp_data = ACK;
        													flop_resp = 1;
		    													send_resp = 1;
																	nstate = CMD_DISPATCH;
      																end
													else begin
	 																ss = 3'b000;	                  // select Trigger digital pot (in AFE) on SPI bus
																	nstate = SET_TRIG2;
																end
	 											end

////////////////////////////////////////////////////////////////////////////////////////////////////////////////
/////////////////////////////wait state for writing to the EEPROM//////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////////////////////////////
 					WRT_EEP2 : begin
											if(SPI_done) begin
        														clr_cmd_rdy = 1;
        														resp_data = ACK;
        														flop_resp = 1;
		    														send_resp = 1;
																		nstate = CMD_DISPATCH;
																		end
											else begin
	 																	ss = 3'b100;	                    // select EEPROM on SPI bus
																		nstate = WRT_EEP2;
			 
														end
											 end

//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////SPI sends junk value initially ,once SPI_done is high it goes to the next read state ie RD_EEP3/////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
 					RD_EEP2  : begin
											if (SPI_done) begin
																		nstate = RD_EEP3;
																		wrt_SPI = 1;
																		ss = 3'b100;
																		end
											else begin
		 																ss = 3'b100;	                           // select EEPROM on SPI bus
																		nstate = RD_EEP2;
 														end
										 end

//////////////////////////////////////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////  UART gets the EEP_data and then once the transaction is over it goes back//
/////////////////////////////////////  to CMD_DISPATCH  //////////////////////////////////////////////////////////
 				  RD_EEP3 : begin
										  if (SPI_done_ff && SPI_done) begin
    															clr_cmd_rdy = 1;
    															flop_resp = 1;
																	nstate = CMD_DISPATCH;
																	resp_data = EEP_data;
																	send_resp = 1;
	 																  end
										  else begin
																	ss = 3'b100; 
																	nstate = RD_EEP3;
													end
										   end

////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////defualt///////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////
 default  : begin
	 SPI_data = 16'h0000;
	 ss = 3'b000;
	 wrt_SPI = 0;
	 send_resp = 0;
	 clr_cmd_rdy = 0;
	 resp_data = 8'hA5;
	 capture_ch1_gain = 0;
	 capture_ch2_gain = 0;
	 capture_ch3_gain = 0;
	 flop_offset = 0;
   flop_resp = 0;
	 flop_gain = 0;
   strt_addrcnt = 0;
   en_addrcnt = 0;
   set_channel = 0;
   set_dec=0;
 	 set_trig_cfg=0;
	 set_pos=0;
	 set_sum = 0;
   dump_en = 0;
	 nstate = CMD_DISPATCH;
	 					
           end
endcase
end

endmodule
